-------------------------------------------------------------------------------
-- Title      : 
-- Project    : 
-------------------------------------------------------------------------------
-- File       : 
-- Last update: 
-- Platform   : 
-------------------------------------------------------------------------------
-- Description:

--
-- Jos� Manuel Fern�ndez Carrillo.
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity my_entity is
	generic (
		
	);
	port(
		clk	: in std_logic;
		areset : in std_logic
		);
end my_entity;
		
architecture rtl of my_entity is

---------------------------------------------------
-- CONSTANTS
---------------------------------------------------


---------------------------------------------------
-- TYPES
---------------------------------------------------


---------------------------------------------------
-- SIGNALS
---------------------------------------------------


---------------------------------------------------
-- COMPONENTS
---------------------------------------------------


begin
										
end rtl;